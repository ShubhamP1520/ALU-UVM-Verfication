`define no_of_transactions 200
`define OP_WIDTH 8
`define CMD_WIDTH 4
`define SHIFT_W 3
`define MAX 255
