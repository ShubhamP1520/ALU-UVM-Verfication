typedef uvm_sequencer#(alu_seq_item) alu_sequencer;
