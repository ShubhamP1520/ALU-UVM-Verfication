package my_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "defines.sv"
  `include "alu_seq_item.sv"
  `include "alu_seq.sv"
  `include "alu_driver.sv"
  `include "alu_monitor.sv"
  `include "alu_sequencer.sv"
  `include "alu_agt.sv"
  `include "alu_scb.sv"
  `include "alu_cov.sv"
  `include "alu_env.sv"
  `include "alu_test.sv"
endpackage
